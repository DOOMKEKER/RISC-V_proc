`timescale 1ns / 10ps
`include "../rtl/defines.v"

module data_path(
  


);





endmodule
